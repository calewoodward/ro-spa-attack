    Mac OS X            	   2  �     �                                    ATTR     �   �   J                  �   :  com.apple.quarantine    �     com.apple.lastuseddate#PS 0FD0081;6577def7;Firefox;CE445F4B-648F-40FD-9C27-2AB8D00C91D8��we    H�,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         This resource fork intentionally left blank                                                                                                                                                                                                                            ��