    Mac OS X            	   2  �     �                                    ATTR     �   �   �                  �     com.apple.lastuseddate#PS       �   �  "com.apple.LaunchServices.OpenWith    �ee    �uq    bplist00�WversionTpath_bundleidentifier _$/Applications/Visual Studio Code.app_com.microsoft.VSCode/1X                            o                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         This resource fork intentionally left blank                                                                                                                                                                                                                            ��